`ifndef DEFINES_SV
`define DEFINES_SV

`define RESET_ACTIVE_HIGH 1
`define RESET_ACTIVE_LOW 0

`endif  // DEFINES_SV
